application.name = Feedback
application.createdby = Skapad av
application.index = Nöjdhetsindex
application.edit.error = Inmatningsfel

application.error.loginrequired = Du behöver vara inloggad för att komma åt denna sida
application.error.noauthority = Du har inte behörighet att se denna sida eller utföra operationen
application.error.pollnotfound = Kan inte hitta undersökning med id: {0}

model.consultant = Konsult
model.consultant.firstname = Förnamn
model.consultant.lastname = Efternamn
model.consultant.email = Epost
model.consultant.phone = Telefon
model.consultant.administrator = Administratör
model.consultant.password = Lösenord
model.customer = Kund
model.assignment = Uppdrag
model.poll = Undersökning
model.poll.contactperson = Kontaktperson
model.poll.ongoing = Pågår
model.poll.closed = Avslutad

navigation.polls = Undersökningar
navigation.input = Inmatning
navigation.consultants = Konsulter
navigation.mypage = Min sida
navigation.logout = Logga ut
navigation.login = Logga in
navigation.home = Hem
navigation.new = Ny
navigation.edit = Redigera
navigation.reset = Nollställ
navigation.save = Spara
navigation.cancel = Avbryt
navigation.score = Sätt betyg
navigation.delete = Ta bort

error.pagenotfound = Sidan saknas
error.nopermission = Behörighet saknas
error.heading = Hoppsan!
error.login = Felaktig epostadress eller lösenord.

index.heading = Välkommen till Feedback
index.description = Feedback är en tjänst där kunder kan ge återkoppling till Crisp-konsulter.
index.guidance = Om du är kund till Crisp skall du ha fått en direktlänk för att ge återkoppling, annars be din konsult om denna.

login.email = Epost
login.password = Lösenord

polls.poll=Nöjdhetsundersökning
metrics.create.question = Hur nöjd är du med Crisp och {0} idag?
metrics.create.superhappy = supernöjd
metrics.create.select = Välj en siffra!
metrics.create.higherscore = Vad skulle få dig att sätta en högre siffra? (frivilligt)
metrics.create.name = Vad heter du? (frivilligt)
metrics.create.closedpoll = Den här undersökningen är avslutad

polls.edit.title = Redigera undersökning
polls.edit.noneselected = Ingen vald
polls.edit.error.customer = Fyll i vem kunden är
polls.edit.error.contactperson = Fyll i en kontaktperson
polls.edit.error.assignment = Fyll i en uppdragsbeskrivning
polls.edit.error.consultant = Välj den konsult som har uppdraget
polls.edit.error.createunauthorized = Du har inte behörighet att skapa undersökningar för användaren {0}
polls.edit.error.editunauthorized = Du har inte behörighet att redigera undersökningar för användaren {0}

polls.show.title = Nöjdhetsindex
polls.show.score = Betyg
polls.show.nodata = Inga data än så länge

users.edit.title = Redigera konsulter
users.edit.error.firstname = Fyll i ett förnamn
users.edit.error.lastname = Fyll i ett efternamn
users.edit.error.email = Fyll i en korrekt epostadress
users.edit.error.phone = Ogiltigt telefonnummer
users.edit.error.password = Du måste ange ett lösenord, minst 8 tecken
users.edit.error.notuniqueemail = Epostadressen används av någon annan

users.delete.title = Vill du ta bort konsulten?
users.delete.info = Du håller på att ta bort konsulten {0}.
users.delete.confirm = Vill du fortsätta?
